module datoentity ( 
	a,
	b,
	c,
	d,
	sel,
	salida
	) ;

input [1:0] a;
input [1:0] b;
input [1:0] c;
input [1:0] d;
input [1:0] sel;
inout [6:0] salida;
