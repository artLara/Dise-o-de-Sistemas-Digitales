module p1 ( 
	a,
	b,
	c,
	d,
	sel,
	ref,
	salida
	) ;

input [1:0] a;
input [1:0] b;
input [1:0] c;
input [1:0] d;
input [1:0] sel;
input [1:0] ref;
inout [3:0] salida;
