module datoentity ( 
	ref,
	salida
	) ;

input [1:0] ref;
inout [6:0] salida;
